rsqrt_LUT_inst : rsqrt_LUT 
PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
