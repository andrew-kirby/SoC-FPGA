library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity compute_y0 is

end entity compute_y0;

architecture compute_y0_arch of compute_y0 is

end architecture;